library verilog;
use verilog.vl_types.all;
entity rf_testbench is
end rf_testbench;
