library verilog;
use verilog.vl_types.all;
entity dp_testbench is
end dp_testbench;
